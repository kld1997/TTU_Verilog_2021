parameter PRESS_CLEAR = 5'b11111;
parameter PRESS_ZERO = 5'b10000;
parameter PRESS_ONE = 5'b10001;
parameter PRESS_TWO = 5'b10010;
parameter PRESS_THREE = 5'b10011;
parameter PRESS_FOUR = 5'b10100;
parameter PRESS_FIVE = 5'b10101;
parameter PRESS_SIX = 5'b10110;
parameter PRESS_SEVEN = 5'b10111;
parameter PRESS_EIGHT = 5'b11000;
parameter PRESS_NINE = 5'b11001;
parameter PRESS_NOTHING = 5'b01111;

parameter INSERT_NICKEL = 8'b10000101;
parameter INSERT_DIME = 8'b10001010;
parameter INSERT_QUARTER = 8'b10011001;
parameter INSERT_HALFDOLLAR = 8'b10110010;
parameter INSERT_DOLLAR = 8'b11100100;
parameter INSERT_NOTHING = 8'b00000000;